-- megafunction wizard: %LPM_DIVIDE%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: LPM_DIVIDE 

-- ============================================================
-- File Name: SA1DIV.vhd
-- Megafunction Name(s):
--          LPM_DIVIDE
--
-- Simulation Library Files(s):
--          lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.1.4 Build 182 03/12/2014 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2014 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


library ieee;
use ieee.std_logic_1164.all;

library lpm;
use lpm.all;

entity SA1DIV is
  port
    (
      clock    : in  std_logic;
      denom    : in  std_logic_vector (15 downto 0);
      numer    : in  std_logic_vector (15 downto 0);
      quotient : out std_logic_vector (15 downto 0);
      remain   : out std_logic_vector (15 downto 0)
      );
end SA1DIV;


architecture SYN of sa1div is

  signal sub_wire0 : std_logic_vector (15 downto 0);
  signal sub_wire1 : std_logic_vector (15 downto 0);



  component lpm_divide
    generic (
      lpm_drepresentation : string;
      lpm_hint            : string;
      lpm_nrepresentation : string;
      lpm_pipeline        : natural;
      lpm_type            : string;
      lpm_widthd          : natural;
      lpm_widthn          : natural
      );
    port (
      clock    : in  std_logic;
      remain   : out std_logic_vector (15 downto 0);
      denom    : in  std_logic_vector (15 downto 0);
      numer    : in  std_logic_vector (15 downto 0);
      quotient : out std_logic_vector (15 downto 0)
      );
  end component;

begin
  remain   <= sub_wire0(15 downto 0);
  quotient <= sub_wire1(15 downto 0);

  LPM_DIVIDE_component : LPM_DIVIDE
    generic map (
      lpm_drepresentation => "UNSIGNED",
      lpm_hint            => "LPM_REMAINDERPOSITIVE=TRUE",
      lpm_nrepresentation => "SIGNED",
      lpm_pipeline        => 6,
      lpm_type            => "LPM_DIVIDE",
      lpm_widthd          => 16,
      lpm_widthn          => 16
      )
    port map (
      clock    => clock,
      denom    => denom,
      numer    => numer,
      remain   => sub_wire0,
      quotient => sub_wire1
      );



end SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone III"
-- Retrieval info: PRIVATE: PRIVATE_LPM_REMAINDERPOSITIVE STRING "TRUE"
-- Retrieval info: PRIVATE: PRIVATE_MAXIMIZE_SPEED NUMERIC "-1"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: USING_PIPELINE NUMERIC "1"
-- Retrieval info: PRIVATE: VERSION_NUMBER NUMERIC "2"
-- Retrieval info: PRIVATE: new_diagram STRING "1"
-- Retrieval info: LIBRARY: lpm lpm.lpm_components.all
-- Retrieval info: CONSTANT: LPM_DREPRESENTATION STRING "UNSIGNED"
-- Retrieval info: CONSTANT: LPM_HINT STRING "LPM_REMAINDERPOSITIVE=TRUE"
-- Retrieval info: CONSTANT: LPM_NREPRESENTATION STRING "SIGNED"
-- Retrieval info: CONSTANT: LPM_PIPELINE NUMERIC "6"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_DIVIDE"
-- Retrieval info: CONSTANT: LPM_WIDTHD NUMERIC "16"
-- Retrieval info: CONSTANT: LPM_WIDTHN NUMERIC "16"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: USED_PORT: denom 0 0 16 0 INPUT NODEFVAL "denom[15..0]"
-- Retrieval info: USED_PORT: numer 0 0 16 0 INPUT NODEFVAL "numer[15..0]"
-- Retrieval info: USED_PORT: quotient 0 0 16 0 OUTPUT NODEFVAL "quotient[15..0]"
-- Retrieval info: USED_PORT: remain 0 0 16 0 OUTPUT NODEFVAL "remain[15..0]"
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: CONNECT: @denom 0 0 16 0 denom 0 0 16 0
-- Retrieval info: CONNECT: @numer 0 0 16 0 numer 0 0 16 0
-- Retrieval info: CONNECT: quotient 0 0 16 0 @quotient 0 0 16 0
-- Retrieval info: CONNECT: remain 0 0 16 0 @remain 0 0 16 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL SA1DIV.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL SA1DIV.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL SA1DIV.cmp FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL SA1DIV.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL SA1DIV_inst.vhd FALSE
-- Retrieval info: LIB_FILE: lpm
